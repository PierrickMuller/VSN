
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1_1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
nyIOaahx/faRQ13ZqwKqvm76SFW4YontKM9Lk/fvFRaVzCHgajKcU+tvMf3TBPWx
3BnsXoQ435sYKHgKjvJnA1UW8dAHyF9rMYbNLkNJnDO3DRS11LMzYj/grsR7gQWL
oyJUB6Z/uo02KzwfbmikusdU7dTuwhUW0WIEGi2tLNzzMtpEJmgPo+FtmWuA7x05
1uYAHHgYjtucgDg7L96q7PAWo9359Dk7qF3r/aS7iPrfX/QupKWH9f8QUhDTF5aF
rVeVgaQ4SqYmIPtIZgzrTcgfJRLKMKb/7lLhKylP2TGmPNpFDkp9Cy97MyxNrtsD
2fIfHQ7sTAuxoOmdyrUyUQ==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 2160 )
`protect data_block
ex9x1jQS81Xcdn3XyKApvPQs6QoNhP59YPEI7m2msWNbNZFBo9wBGPv7ybWtcsNU
xA+J1kMF69it/Ri3IG4I9ZvYsa0s5xzWuchio4waaMa38Lf1LZo+SyeJ+/LUyqNt
fEr+NTATvNovMijlHT9MMhhSdHNwQGw1F7I0aab4hiZTzsC2ofExn/F9pusfAbtq
aFjmg+oQNrLgwpSRV4yoFl/fUW4g3jFmlvgDdw0hVW0mANcZsL2tv+ndsAnGFCxy
55j/2udtiB3p8r2oi46MTZSiylwUteQwLEpCxVi5CdLmRcTuDmtELIM63gI+w0kX
HAz6EgAqBHzkBeG3IrGhJaj0wK3TW+maxEjjYeIvc/E3hTKGzw7gd9P1InoA3Bz2
DVgv0uzxmShHXj0ppBfvhZgQRsDAmTOAOx7dbHvjsA8pbWjt7nhkYY4+oJCXq+mH
obdoRwCRmtMlopz1kBoCoXb6gJpJhP9DJmBkp6yAWt9iN7aM4ppjheixjmmfNlBf
iTA3g7TOpn4QXvSP5uuwcycvsINsEIIDv/5P8HQxfKpNvGEoGflW7IetuUF5Pl4D
zjepNRugkFnCtRiNpF0ZBd6oOCcEis3x5bqhacCNsHaTdM+SbKitxm633BLcVLwW
Gu9nyX/XzGa/ECYRrItsxkZWB6S1CbtvRtu+CFsZJ2iCL4OYboWVK7oai5uuEgXg
zZ02TUOBro6fFyJXGqD5IQxGj05NBBldELBMMsly3gRoc011eff/0UQiCeqQ0xgv
HJKULh87r+OlL1KZr12VgmQXmYZlWP8GNc8CUcfQcRv17XwUi9H+E+WytWu02C+e
esgHZufdjSlizsGv9rdj9Pz1LuHKsIVbsxXt8uCcTDRLeGBZgPnWNZDoRHLIRVPe
cGSDVf00ExhSjlBwfxxXq+FMGg33UtmM+joNWuzZQSjGWHY8RcnGCSSzq4XMTlT7
iEot8mhZRxe/s4A+nKLXDrFQkEkiK4yRHKa+Imrm4w5sQfFh0y/ovmL4o0ijBOwm
IdglSmtGTvO+imaBDRwWDhsSqjlnkBf3blIF8fQKjl410TVo3KAXnlHc1kXL0+Ms
jJOJc4qLbD5Ik5IzC56mU5d8+6aAsf44Gn52N97521vKWh6RKEqWSpggYITPxQmK
HWNH5WefVqjr3ZL2Rm/cgCVXaW6TdG/IjtBdyr4tIxeOrNAVygoXN8vUtiIgJQi+
f7FS8V500+ANMs8NPj8y7uX59sSTJQJZxThWwmAUAVTtv+ZFUR+E0raroOS/fFYS
ynov+2Jlsa7qpWMq2bOawLRdEVjZ92jmsKiXO/Dj5E//RIe88KMIuPM4zT5qdOyV
T6YMK3vUJtaWGPDs2kpc3631cs9iRXahJN2EUjT14wZtcr3h2GeE12nuuQjxfCGZ
domqFs5etKCSYL1egt2kb8ZdWW1QzQ9Iyi2lwsH64MHoZLjlrL5tl6IGB3jxcgUt
QdLQ9Q2lBasL5Ytywl2qp0I7Y4e8k9Dc0seJ5bjGrRceU2EFVLQrrqlvPjfy7of4
yoVeWl0R6lym1B62G2k/RmjbyGTPLDURXOD+M/yf0siXwoSv+eGm6MPfpY8P6G+G
dR1ltJeZgsTelR1FubTFwDinll03wjzA7p+rgmSBJdLEZ16Pc5Gx+dADOivINVJG
KD3E5g0x/7tpeV36yxJ7SziL6vxIe2IWVEt3kqxic0KOEjZ5IxxCScUOvkZ6bRZn
ZEIhXTKfZRBnbYSTw2bsGue2T4zsL4engh7vasRAx7iAl0O4niTH7wMQor4wQkp0
8C+xQegumuLbnQcJNZY1lpjRCTjeYR/w6mCnoHtlzGLyaRVNTrYh36hbFeoCBmeU
wnPi+dkgSeyWjuwGiO0nl1Qxtlcs/o4Qb6U9r+/cLIcyKDt34h2qLRTZTiqRe65Z
WT/mAn/sziVzGt9lB8uy3zLbXOtDwHPT6W/yqQt5Xt4gi2guEWQ1hsYgZw66FUAZ
ApBrEmseKfvhxSJ5Bj6DGnx9GyoBX+1W9bMrmeWbWLW06vCtbKCsurhKm9jn0raP
99Io2A6reGeURg72/LDz//0DPrEKsv9n/lDcb4r6J66zeRZfkBXEwoWdpavKv2x+
nnmUDvy8AfCNuP6BRDQQy4yJif5VDbbwi3nUGs9iqqq6y2fSyioNhRajhLLs9p9Y
hiFEdG1SUMs9KkNwdi6wj01QTA+ZmeI2G5bJlNS3xMLfkNQPcqc0UgKgwgpSJIMX
a0SxsiRlWgTpUzMt480B+qjeVOP5J8IvsGc7FbkJAhNl+TmlF3NEVDr0GjPfLvmw
gt3p+rK8P4woh4QEvkeIp5HpQubMhbsNNynbIIST6aqutfbE72qKXryEowtqVeDa
qbDmQrdP2r9Q6zCFBH8Jv+nUH3Elf8pvKo9y3Q7CYZCDT0IDUYnH4o49/NTPKWAi
O9rgMIgOUmlkOHzGiFl8uXrCaiw7A5PJ/q9Wfkx3DPAH50Np/AIjntP75MnnM+0z
I9gg5UmH7OAqB/wfODGrDz8oDJ0mIG2UeDe2FStbXgV0xZcnhnpsG56FTonzFvqO
SKRpFrnD2/E95eXE15qOfUsnuwsKrkS3tHN/dB+3R97UF9XxpoJBifx47GssSrvv
Tc+7Fm1SYXLQlVZb5oJPF0AOi8PIpEDsSeQNZcDerATiUIqiZWXnKLfGq6CUkEQx
UZdyWGJg4VQO6RTb63Gaet+wJd6VbFF4d6OsN0m4QZUCU+JSMV6+GMv88GsLlUNt
qG6bEKDXRLPaLSXYpt2xFKe5C97gg8KvZSNrp65MuYcp4hl2nZiH0hm7JgF2wSjD
p2tr0sxCBQdDl7p4g2Rae2NA8G/qNyU3pecW7l1NpNEkxL9o+36FJ37GONDp891a
`protect end_protected