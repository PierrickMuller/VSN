
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1_1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
VcdyGU7ZmWnXgqCLcjfcDcCOAuXhu7yXLboaCzOJHKT367J/bwiP/UuHQB+EajKf
5FgV5dlMRKaCLHbysNuf26d6woFy5Zm1tKbpefEDlD4wURUy7z8GImxlTFMmSbpK
4cFBxtNn5UHfEpoWvW9TukzrmWzD515+UCzND7+UJsosrrTzTovMnG6PAp8YiUFQ
ZJTv5DT+wN5kkaMLV04R69D7uSjWC3GjLM3vg4CB6+By67XpVGETcgW11jo5tYCY
rDdWwVq6kqZCULC2tFR+CDcwFXpN2q4pkZNvYt16yrImQZIKmOeBIiAajmTt5TdC
kCflTDQ3W3Z6jwjSVGlJMg==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5440 )
`protect data_block
GsjZUbij0rvb4RimWoWf2OXMOQTG/m57ZjmHrI4/TFeNWzXnBt7+hd+tPi/SuEz/
6BZIG3430ZAGiyPLJyKTtAC8y73+gpAnOxqfCMqXB3xBWAvSuAaI66krTRMr6S+s
dS5VcwyA783+IdyvyCbbzyTfaP5LC8B5hXOYSudAr1jPYteVh95z6jaVuNQPOrdR
Csksez7SrSlSSIONoCBn1HpHkNXZVESU2W5SOOqPHgfc1FsfG9l8RU5c98njXuV8
gXZDbFIo2AehCpWuX+5UC/6SExiHGdEoPidaJksIoCRBb2xw07MDNB7AsENC2RVq
+mMpr8Cr6cM34P/0moQ9DG10SpCbpFuaxSNb4+YkAUykG23P63GUzMW2cdp5IqX1
oxjaTIKKR0QqKvf8w/DT3UZAIJrW6zeD+WqjABS+LBQIHKXalvjj51wCBxEotgn6
pR6lQArXcthrmdjGskbjUo36hJbBpyQyh2bS6Qry0+2qhf7QJlCdXiWSVKJN/D5i
wKUNtTRai8T92sqwDNd86+VLdtp/h7aAAak9xNBf4iPCcL7enZU1AsNhhjhudYj3
9tquP2w8iuCUvdPzedddElgQ8MHCNvs4XruKji/13UyiDP+Lw7oYetAtkv0a4W/H
P05f2NPd1MQu1oyOTqkmJPuRJ5/Oj+TsIso25nrBU2PTctkY6adoPYGRGaQmmu+I
NQMcyHSLjgOsW2t+u8e+Se4ED3I+frvXBjwAB+1oG4ZAWeRRYASFDWxBeUo2wkU2
a3mwj5MJmPrZznW/4WT9+0NW22yCrImX98nKNNYbMDzztiEA6IgiYXNHjjGzwXOA
mtZtzskrdz0+D3AdE54chHVMUdbpMwfcw7+pkEXFoGcQfTKuAAHqd1f7G2dp3Cnq
oRl0mndJGVqUzOxcb+4QYzH47U/ekK2eCkVmoUaoFvgWU0KPxPrZ+51/wfnjoIgB
nV4MiwJX7YPlh7A/s0efoSb5cpr4on+AgveXA4OIQvkBZqB+6FXKkw3iLn3niUBk
jHU9LXNMsKlHQsikVwBeXFev4SorTZhQ9681HPlF69KPu/ldNDOWvy0D2kglxKZF
QkeNesCcD5jNgR/xeEleWy60uHXLKkga8aYI/5p8OV7jHa8/JYa9WS7VV9YTjLOd
jdjwJTTE2vjHMyWq7Z5O8XRl8Hg+zSzztkn02uZbwE8lXpYPLbi0tp5uTMMfjRmM
w/mX/32cGaBsSORIgroijL6ktoLkEfNWdHKFx92ALCTiDJTSzQ/LqCB5EbJBjG83
DP8OJqqe0W+I7Leja5gj/tQFlLn/z8vRQGqKd+mz/qHHb74FnbPGQjA0XTqpQSs+
o27gPNnTOtPxGEtjJDtdp2zj8ULXWe6XC0KxsiNB39A0NXYln2wX/i4jxFgwI7rQ
nakZnj/VoQ7eCJxDbPne/fXauz45NrKwNtRq5Ef6+T6VYxETxNpO8V+PM91ZAKFw
S+4V683zFIBpl//lpDhLiwEKTmDC4BeX4sAB4NNe38mc8bLkq3vkGmDthTl1N7bt
wvYdKowpv6RGUTqOIqXtXzCF7zLaoMa89aUDOERijkuQ9NoCSuo9Bpe4t/OEs/o8
sFtuq8K/gouCCOAeS958tJ22wijvOSOqJziB3yV6MloP+4NqL2G3qKi3grwnQcFQ
QRRg7WtjShFyw8rWYh4kZA842/UPSvqjx+UqWfc/DuYtto/lxp74a6EK/tKuIW5Z
MkXyCz9uEIG90K5Z0qw9puHm58Xg3kcoeEeiTSlB48hCUZKEsq5k23Zsb7lQHdNb
FgoEIRIXi64IsAINHdf0j5xLefakeZJzvH+xs5QSH0ylRqyKxzqgXJmCCJx7dGd3
RK7cktzXjnydfZfBMR2AKiI75aT/lw3Klafm9rLO4JzA05JxsrCPPROZ3xH7nXQN
EwMQG25UsZ4U7Pac3O4z/pyc3Td0rYH1jGSrJkKkfb4t/+viP2KngFs4lCqMzvYL
70hztrlDecV9O5vQnrlNK7Oj80x57gWj68sPu2hMvbtRrqM9Pv3w50Oi4u41jm8p
Mn/t71DLCfcqS8uhF+2HQon48Fwrm3AbtXNsZQ5Lc2squk5Mf2zlofUYJTMoXPDi
cdl15PX0c0F7LzO8Q1vKDApTtLaNfWg4GVsqC4aFB3eHo40WCnCZSZ05Dq65NURo
SVWFXo3gcUwRfkADw3qgIb32jL4klku+hfaX69ERN+2WvAXZc5Nhis3OYir1Xe2C
rMXrALj2W7EtEEh64ZU+PC3lrh2fbEEjNtOThNlGAa1rhkLEWsNeShE1EEUrtFcG
SnZvq9KZgILJZ44/Ul+jzuwGsuflcPIjYLAe8x1GMJDn8fGlaiyg5UC3h3ygayxW
zfQkj98hD4fPFXt3+Z+4SaCoqF2dZv6+tEdzh4uL0jJlU/xVMkktuRfI0Jnm69Ni
R2m2yaO+74NTTk12M5KsBH2YdQcRWSrLtb0WbyVMK9tN3Wi+PzH9pxLAHxgUl0fT
8JaUYhq9soXiVzYh8YN36mkpaCKJzs+8+ZJQqDIuGusu5T1jdzY016pPZNWPE1iU
IIaUoA5yUkmIwv5EFk9r5Bs6UWrGDltMHbuoLetfGGE1YWLwRkwmuMbxCAjSH9OT
FUHqG8l4NVJK8KI3ujWCPr6dRe56/j2HeQ2PNWxOKpTBJ28J6vtIeLQLyu+7P79d
+4tqZ15kCrKS5dHz3TR/QBtdCGwAbhupnGSTnL4opmoq9eQkFHu3mNzWvYC3YajF
Tkax3T3ToOQE1P8KXR8jwun4OJe7RnB0ymeud6JRuIXnNeIl1ePF/3ufkziLN/jZ
OvLzs7cuocv16/dwLlOBEEA7IQqGdavuPETjvCHOygcyFAwsz1Jm4zUjQvCbQq3q
J/IImjFJo+KPS8mpDorZJyNXaLms7yg1a+SJwBLythvxU0FHXZZzdPlcRbyT96kj
V28ToMt5uiXe7Vq4HKdAN13L8YCD9MJ/ZAUanxHGbAkyr3Ezu9Mp3OAUQ4hJVUDd
50KzM6/tTXd1aAFKXpIa4RmZBjpWXQ/kaMnjqM2vh/XA4MN1H4b0F95LsbAMoY74
hwKTlaYsFv8AIt5Z1kf+EfPyAe/+Um1mQE/ru8yGeKNb2wj+GxdRi1lrksoou26I
M7EUJ9Pg9RZK5ptConevKDM4v53H3lG0ryDXadeRsBZWJwgUHoURbGHAttOXEctB
ucPcHOxly805flb2nLuA23Mu+8AwFq6Tpnv1Q869kBAeF3ttba/DPVKYqxDVt1EP
jFDvkeuVM9v8DaJOIA2dobWtl3wQQZeaThplN4/V7L2rMl574i7+S7fLfR/S4bVr
filKd8ujkHufaM8nzvf37jtPIQuFE92y4+C5ANLFKa+viwn+UmGr3u9Va340mB8H
9jg6Yx/4+JtCC71dkHwmKKyqiGXvA9K8DOVayFbPs1hsKthuNFSjHGlTkj0kzI5S
wFg22hnSZkquVwIS53Xd8AWuO2Xqu4ZadMPFcDcG7F7c0QalEBqWkGMZ+HW/bRdp
S4CuIUqqVAFoVN6wyLKoxlMPI/v+vTT9N/ZXwDVpAlvRBcczRo5VeMuP3/zT8F8l
diCvihZ2//gCQS876w7ci2F75dFLl+c2eXoMAppram3FRhITXkzDX4XWRW9VAWBF
AfAzB4P7o+UArmlc00Pz40/iYQMRYw7YQ1e7MlIj0HJdVErq37mKIWkCexQQnloV
pXQFRWwhNObC8q48MsfhqMy3s1GrkWhJVvJTuuZK7C1JPxjKH2EkU/nL6v4x5dCk
SeKTlplbpr819a9hSoWMc+Ku//sFH9LrM4Ki1Ax9PGLFT66cI/5BvRK3pA8Tfhi9
9t59czn1FCQqskkt+QLbPvRkUaYaQpHV1jQGR1F1+hfA8UlR6etABIlO2Kr8uDMh
27vUk4jh2oOe5elqq4nO1eJMqKQvr0l+3c38TNdHpJLTS5R19JMyZxUrtgTiAuXn
4HFleNPukJJ0SpP47cBdfAlOf+KbEpbWJtLbf2EH/lZ7AlqmWuwcYOfMKyZIUCx1
P4L1LUGUuWr86v+LyyrYmaqLjT4+XhyboB3VxzYRyoz0OyJ6VvRShfM+jkaudlbL
+BQsn8/TC8QDaGkcC7+alx85arpiujU/wVcq+LzlA3FL8cURpEFXd+lYG2L++SRZ
b+Kobvv4XP0NaGqM6H/W6jUetkNOOvnwPcyxmFckeMBTWApXib5UdDA6bq9lwpjW
l1v6OlcYtbNCjJWuVtd/FYxiR38LxVfGxnMjYMFtmy2pZUb8AbCadPdIHJCLvR+i
t+84qEFwT2mw/mFDlVTRVq5I6lNKDRBnLaVkSk/G0JKKkxlERUvSvGERjtIS1dG2
9H/xIqfxd4w7ZaPEutEDV62Pj2Nx7ouPRJ9BuBzrKysQul5U8F4b0qtTxJkXMA/e
jdS/f5YLYv137dezZusfEIV0ES+L6XUmTxm61ZGA7o9rFJwUY1S04BaNDigLTw3w
2eltik233R/Ca20oxrZdG81cQJ3IFmM3wcETXYvIsNeIEv//Io9Ik9Y/fQkhPRQc
1s/8lmT/SijAfLYj0f9qo16HveB6A1OoJsOHRl9taC4HTg1wiCsVCOI4Q7fcXUQN
E64MJup1Mb7fZ1N3P/mPw1rzGJ7+bPt+I9nM9GWlM6QfKA4hiFFhgXWWt7mCF0ud
fAmIt/wfvdMqmGk33NMHheuqS9mnadypwI+9yUBkuMAXHRDNy0AwKLS4tceUSmzJ
1ckLYMhqk9GdxknRyMfWiQhOAVsAk1KOMgfU4Dv1EFgXhHPBWUk+R0c+xgL1Hias
biLDld3Rb/OYHmlfktKXwaBwzvC5K4zEGjlSYqXYSFULT+icozclRvclzYAvDJIi
3HB9GwFm4AFzOm4m3pEUEbVHX3PyAaCBFF4alyTqR+89QRXGlu9tRcYUYrNToJYr
v1lKmhOqjGj3sgQ3czSKmuj8D/Ea6NZHviuz60m/rUpDSgSwZLVohr1+tXbXMiDw
fydq1iQn9FPFLAZvOcyxfd1D7g0jAO1ttQbaKmeS1cqhwMYTE86LvagGCb7KOXJu
kZP4s2a9oRXXg3aWBY8GfbNThATPbfgWZGMU8ORC9fzGux1Ze/iZNYe0dtJAPiQk
MtV0uM3ZW0377GetX91tOXRqt/cF13aQKthlyB5m3pCyhQ0GpZHwG3HdzGvdwJBd
r1Lv+soOX4Yeb89AGloFybT/jWpzLw/SUGjOxBFgAKvgx4eKJZv2uQamnpMfQup7
RdXh9lPhMNjwFnSx/QZDCkjKwMGbghZe+Z/gTlOn9R9YEbe3kQzRGk2rUguNoMaR
VDnZYhAml2Nq1eLG2FG1gl221xz80k6EK9fA1UGiZbKuu7bkLf5nA7sIRJ4bbDRB
XxjbuHHaVpJ2afUCFFSXpUQk4JodugZ5IeKE7cIWWIRMjWWnfS19PeaRAaEwKi9u
VwRIuBsUXfCGnP1h56lqOto0b/cI47RyupDB3cwyiDNqQEhVVx0KAJIWKWlkDcmW
HP2ls0FL4P7BeWpfPVGRFWsUxhlQALwEaGPpV7CguyOu6ZH9MYRRSiiizHcr31w5
bvi4c49/5ZeqPeDSjmOEdPLI1FiWw9RBEl+MhxLcLesd6BU/tRMNZKhznq1u2tkw
niF17odJthctV40GMKxUad2SVbYWup3b/cs/COIfns5BK9h3J4kV9sYPNiHH83ZN
DHRaoTr1WQ4GAeNTctnfK/6hVDhYMk1Uqkf4bdO30SyUa2NUopj0VYQ6+9cPH1xL
Dwv86Yd1tws9JFToT2YLaG4Xgu68tcBJlm4q2rndzNqDfD7vZfgGIelF9y8fk1L6
YF53sWLlmTgelUi7nEe6Tj6rmbeXnoqXH8PUAbyHkc98TLvB41vw/6882UbdqnMs
m2RCHL0xN0c0XQyZ+0IVCd8mZuNXkMs6x+KSN3sXz2SeCuk2BHQXO+3ZKsHJ0VQe
G94PFthGauaiuBqqOcmUXMzRwSVN+AIHgxMrFSYeQpvNfriCzi0iWErzH6a+6K9R
o/09D92fax7/TUsGunm2LzPiEzj9EetuXVRiuZC8Ri0hJjzZty/fXPkvIYtsIssE
cE1fKdN3gH9NRrwlocfFZ28ezQx/Pa8UxqbCnfCLocgwBTc0P7aRvq5W/dcm6z77
25NgDrvoVQg/q02mA73y3hE0THuok7xVo2IwqTrIYS7KRPhC0p7+FB8CrRcEZzol
cm6BNwy1W93mYkSFel6kg2vNPpA0gbx68dQ2z1abzXtWZgaQ50UIh8gqYtJ9JVmZ
SGYrBulkZe50+An1y4Cdmfh5QX95kx06R1X5pOP5ScxIkexHIjMyecV8dORCFUtO
+m0E4dA+s/yM3/g1Y8RgiVnY298a84NHUsIB3VkTy0x2QSM+hBuFUTILz03lj5Z5
BRMpfPgClGxQGJX0jH4m5m8Cht0jQy24APt/mtBo2Mj14UTE5i8e2EB1WRm+NLd5
MgtLO+BfWeDqEnm9md+uBOy+2Cm1KTkzRUClaQdR2H/S0PSfVqztS760S4LVbjUJ
YDpzAHm56hSD0ufcZyUpyjpUwHcMC8L1VsY7uvlRytBXMLs15YV7kJfCUIAPPAWd
HL103JCZSdLA30B4XRpSLLsVo1LAWQKNvmmBmBQ38B9OTva+z6EzI+FrVnXxox5Z
anN/rXEDQ1RBA0qk/owz7emvaWfEFtyiNVGIaKJ/4uYRQrxcaOQ+1CLIjElFW2iy
zMUtmOFMKCrzIUY3zLjFWL4J9HH/ZESspjjSq/53vSggUHQDpZcXp/Vl4OUymgFg
WhHTZfI+WoZjafCaQf2sdzQwCu+3/FUzWY/oomaDlLXtyEZXghRcExgQduSNFk9y
2rS5d5z7n3tokkPDCXo7OtxVqeTV15nokGy9tOQIglP4iL1xPIZNJ0hw9PpMA7DC
S+8RCW+p0lmwS2zc84sThpF870I/8e11wXLoYtzHwYHFm8djkjHhUyM1XBs+c3+J
uEqTGajWD5OKIoZ0FtmI9wUXRM/hSOlYMOg4HN+9hwELCJLObun/qBAK9Sxey6gq
knmzBBHBpewvZ7Q/3PLbbn3/G2igzkaS4G7QqltIr/gduaH82T3jWQRdFEK6hVIq
Sdnm0mE1K8QSOTfGPKcOGnBMLKY24hDl7yD3wEuC6wsm7uPc7lQm9EqTcajHJ8+I
zlhf67Bbf5tDK5jClTkV859fGEzY1LEthaCkk1Qj8BZH1FT/QUKy0iARHsMkXtBT
S2s5VIeZFhDn2glC4ost6A==
`protect end_protected