
context morse_ctx is

    library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

    library morse;
    use morse.morse_emitter_pkg.all;

end context;
