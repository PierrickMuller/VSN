
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "QuestaSim" , encrypt_agent_info = "2020.1_1"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-2"
`protect key_method = "rsa"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 256 )
`protect key_block
Ewv9TuEzDuRsZzKn9Zw0m8ih7OMOrxkORO38SI1miPU7IDQ1gBEzXRKW+9pgOlAz
fkWPdsnUKGNemA8ccTO84TD6bNAoUYBxxcN5kZZFh2uCMD4g7SU0nBFVSPcME3yk
6FErkWog4f460Y7+OkZNRij+KLtJy4cBoBy5dINweVgT7ta8wPW1+ELW6ic7EJaG
Q4nz+MaQ2BFjtj8WSa+1ORYMND7t3jTWJ00CgAXMiAEIozekMz3KuAmOuh7r6h87
bhzhNfPCrmc46N9E8lKBv665crGO8mF2ouP/sSgWI1f+g5+df+AyN350aEd+reG/
mzRHhDDOBzzpSM578vukLQ==
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , line_length = 64 , bytes = 5440 )
`protect data_block
wu5Gp8UMLw5eZnxZcv+PjASjzy0Zc/XWsK7hkTxWSRxPJodXhGiipilBjuBh8i7L
ZTuFbBVCwVyb/Q/OVUy2ELjhe/MVWy3Zf8lOKo2rvE7tDnuEMBpUA6E8kS7Bfebb
NnKbugw+wxNgEKZCnXecVy4yISFP+/ngJs/ZPEFOWqctF/VR360raoIabVJ0fzUf
DIf17/yTwy0lHDDhFr+1TtiPfn60i1tWUpIw7LRxpP19Y1qUx6vgGMbVrKxz2Woe
fkKbZLtIjTtfm4MY2Sv7oRJl3NgJF5AL2qxjEu3w+G9Ezb+RTY6Pqdir4pJtPdT8
Bmr4WckTpSae7w9/3nUZ3pfspXzF8+WiCYEcgdISb30hbhy6/+5EycyNfk0qZn2Z
bSqYV9nUxQrA9LB1t7qICPAmKTWyO6pWHFWQZ9jdhgEmn1+mbjse0bPqbXZfVwEG
j6puqXjOI7Fk+4IHC7Zo5d9QZ4TK14F0bKQRqHt8Rq/01BwfbF6r4TKLHKLMrT4X
6GQOjlm+ZPhAraq+0Rlc9jrLatwtB0rB+HuvnMs9Hw6jD1dVR9ZskjziXMek3H6o
gzn2lr9/JlzQLSl47enoLzXsx/lfJ6zem9RsqCu1BcmCoFAm8UIFHcks/i7y5gvg
aRHngTI85pG5nKl0/ZywGGETA6SvIP5lgxYtOvzRnRQwZXAovxgS7krAAl6zZZ0H
xbRK/UYtTSj5y2sNoKZQcAW6CRZRu7Fu7+gGz+myqcwk5kDFBo3FW+WJjm3nUTud
tu/hTLnLn2/yw+1xuLrMxvvGRnPOqIVFdZcGQzyWAGsjPBycIB12rOpKectVKJnK
qd4FHMjWN5qK4dmEfjGt2FxH6XlPAGxSgSR0pPtL4iHBqqxhXCUGNSJFyoKiwkdM
cd+Nca7KCR52t/VaVr7ys93+VMKxJ9XSmplOuEH36DjxLf8u6y5GEHYSnCT693Wq
vu57FhnD51Dmcka1BDY3vJDhyKbMjKvgwqasQvPXWyKlfzMF10kWNiADmvqVesDE
3WIYn+rmU6fPQggnIqieRFmvGrQqO6xlOkR020TuEAaYffDrcdm1/mqDqt6TnPq5
Po3Zp7zf/TLCj8slAiAAjthLncM3Dio6wkktqjWnuM6MIjXIywB/yyQm57OUgjS4
t0gopqG+ChR4qkp0JqVRdCbxLOcrQ/TXpovZTxrYi2V11qK6Wg3cDYfWwnfnOsBa
5giXk+gqsIEx/JDsWtXCS0yEe/V177WXYCNRoUcQq6VqObBcrR9qOc4lv5vTtZ0Z
wqxm7V0dFPSz68G/gsH4IXYQ7GO0ZCJs2QvQJuO6rgtDVy2zGavfIAS4XHwfRdsZ
yyy/ejr2U/HOxICg1A06sd7IftOVRj6gcTarw2qlYdmu5Alt4EF56BztXtgOMhUo
rze7eAomTgNIzcCnEfBrtTVNxG6Dov/Aj+pV9y/cO7wEL+JzP+68ZOBDeYy7Cdvf
jjQk9eiJP72p8Gn5w8TXuWqthW0IVPtYDaTj5ERTaL+g2eUzcDdU/boXk/cktOzm
U+ufb9JLYa2WBHWEznyC5bqIQUD5ZBCf/1PpUtw63T60R1BQabPLGwJjZR9BkY7i
kSoax6kKaCYnb1atbqmuKGTKVMt36bOmD8ENP8O7tREdo3X9MMMvxVZjXRdg7z96
AyS01f9IlG60YWzfvuoLl3jAv8qC7D+dhGWJ9a0bGbuSN2Iy3BWltfGYuIV0sysp
NWVFCvg/lf1/Oqzbr+SduwP+CbzEdgfFqaFQT3LLV0DSBb4QhxzCa6hC9RXCCTf0
4Rv8sdx1LTLZDigzu9zY6LSso2CuDmXUWp2fS2ysrOZPnELYFLSG8r+odaAdG720
+bRrde/OXDbYJTnHZn2/T06vofMmXZ04rNTJgn0OWoa+syFr6LBHBqarg2XFugOs
aW592UyHco+ll/cZpucilZhwh4B/hSxw3t3zKd9gxhVkDU/pmPb6VuhAwboIf5v4
lFdpY7y0NlzrW/eUnydIRspYI267Y2O37f9pVHlCNlnpq0Gpgz8KxtuMyx/zxSng
oRBF9bmSqsQTV4ftIeX7YtD2n6M57CpH6wroCEfApIX9O5ryVfQ2OuUXgZVz7oqQ
Ez83UbgpF+ZMcBCCHSGYe/aaT+b74q5hAHv/SXztrCVB6qr273at9dyWrmmmO4jw
PZKeg5oykraXPDOl2HnBxf6UhPJ2y2nXTlhQU3S1JVQn4NzG3FkCiTOrCIc4j8pc
9rsuYZNearQvonaNMIHvxddNrecUJ44N4N+w5dZo1wqhLpqBPRb4uPy08Hf/lHFi
m5H6jD7LBnoYn0d0rS5jQZpQdhNgAau31UxowuaL6fPGAusxJYnGwkRTdWmnlLer
jY/arPpwj3hxhTA97q5/TN6VXpdJM5B1Jnp6isIXo3dsma5w6p92ea3B51Bku1+n
f8SmIV/bAu5cdMT8EHkhslZvebH9WsYE0vRlnqFPgLpBHerkz6lIdCxRnetJN/Ud
hCV9++4L56Lq+AG6MaHvIsWIvk3YtD4CVUDkUTomuL0Nx+zeqR/ISmsPe+Z7oMhI
I+IyFDlofU0GhCD9cShebO29Lg+haG1jsliB3tHchBXKj2naxKoYYs06Vs8b3n64
2HbxMDwMHw5o39U5HOY0DOrKktu0QH6+Sb83a6Hkxm72PPLNwb+mBssF4GFJDFa9
GJ3RsvYKfun5RpsibUznurhAtQQouAAlxltDfH2fWe5VvlLHKDNipiWsiW/NGUC1
jvuZYloNI5zlB02aIXn26UP6wBk/xtRERWsRFE7wAsq0FRWDbJ7ErfF5OkVWrQv3
6N4gVOcxdjn0rqpECqXNgkud20shGagJ9yKmY+kjSPGfElryWz9kcf9ba0iL9hcs
npjwZlUDB8fL271FVv2LRFdN1UApDrvWI+u9lfPqdTxDEHXuGxc6KsjZEN92I5hH
K2H7W3mpQCvMaHPBSrhpgwnFOtLm9R+VeYYlySHFNngETwKE0peXiegpvdn+T5PD
bFJY55HKPDvY4/MMMRH1JWgUOUdmON6jn2ObOUomSm4LmbGzeX3B2qsm6PhEV7y7
kuND6h6RnV1N3BXPz6RgSolEH8lOZchdkH2Gaej+NVniMlN9QjLpnYfI+xxdepTy
RFdiQmFajyslntbW+AEj2t2Iwof+UGDiUainvJPd9lNrSGvCCQRxY/k87loLOIjz
nobTnKu+0D5UbCVGbKoWWgvy6adp66PXA5GjhyghWBKkzMkAZC+HtWD2stgxf9EJ
/gitYPMShA5EisDqbgbRJsevXX4ODTvfg8zlQM57Idvanqswtc431M1FW3iOzf8H
hYNNlQ+wEvGgi9klozjhEoXrCk8NO6MNj3dWWMFDBGhl37NsxRl99m3w8r9L8ilu
YKSNPsqh362wwCM718QNAU9vYU4kHGNHsPRUZ5GZdzRkSz+zbgOAXdSBeMaLSuFI
KysBomIWg7d6Du3ELyfYURUHhKvXrRfo33yVlPp3j+3KsMKu6PBtJREFRr195iVH
PfelHMkC07PLTpc6ugtCpCr/D206X1jDkcB7UfutVfZi76B+6yrkuUDkdKa8WbJU
CPXYu0pXFD6IpZ4kOynZFE62a8TgtM+VZxu+uh0ZjLPhn+LxXILFmzO8D7hlQDMQ
r5bs1TIjnbwUpTE0c7g5+1aY3mmW13NxDaQLx71MENKoLRTK/xHNOgnT/NNK4QQW
wDr2mMn9yW2Sag9xEsAl3ZDYppvn21GoP7f4nY8ceyrA0C+O0EqHxnDO8yY6aLRL
DH0GNsN4FbEsPxooWImxe/m4KmUNHewpp7804bXMT543pDPCAk6ojdvr7nISIyZZ
3015PQzU/SJ2D2FKGF8+d+SCAXtLvXWv6ktTXcjsHCR8rDSVF87f+Kv0a7ScHGNP
o6XsaxZyWIF4RH/zwxpClk4+zNcqh9JTbQbLWZ6ESKFOgzZghkKRXL+Zwib1EI/y
F+tYj8bOzqO2ZGDWqZ4CfD4ggQ1J25IR8qaOLziUqNDHkj/bchcdrUHDjl2ft8Sp
1hHz4B/DZTq7oxZ5kVF+9kVzLoYdBmxbjlBdrkgtByA4ZzTBxmmXiPjwV30oHBuj
dDUnrfFOQGXQ4p7pWVE8Yt68fzu6fm0B/rYbj3rB+WrmHSc5t+0NBze1BumQGQ1Z
JGiUr6TWG4qoIX1NDzIp1zipkyZ/5sVkYqwlwj7w6YmBXVFTZSdGROo8j0Q+r9QL
XcTwmjmLepIQXiJ85iGaqeuSjsfPLQRBfN/cFYCy5ScmEpx2eqYt4eITmd2OYlNa
Qv/ujGcYx83+5b6yk6qptpkXF9EJP/0PAUI637GphujbDJLzzNUHRymJNbpSk88W
qSPUfk+QjwLMhBgM0v30erAiQbDxTVGHge1vemYX6QcB6oq4mt69g+XJIyLERxn5
peilPOBFiKVFbGRK/Sx3ydSAtmMUKJhQq8mMCFs5WCbIuYwkkNVCy3ikKuh/jjzu
vE6vWSnj0GlSyJOPq13xglq3C15IgVTSLljULSath95a7jOFAsgYr32DO+z4uXNE
7gE9oOMqpLQuUhVShFbAohSRtu/LdNWS49ukoQBrzI2MZIxk6Y9dhMP/hM4U4dVI
TMR7HHjyNEfaKVB4FwFWksc8amxLjosoJw1eeKWvzti3kLCx1Xuij4CDzoxT+7HC
KwypcNi1x1qcldT9Ynj8Xc0mPGzxi10RCHcvMFx4dibnUsyqYq8noSAVdnFqB95S
JxWS+Cq+HcQATAXsReUO6Gy3JYMlYNiZgJxlOFI8JZ9wa9qU8cQDFNhr8alxOHMf
ZLXM2OBgFDzv2tFLxfoy2YAbHiCI23ER6vctEJVR3jPKReaYHyLy4qt0EGZxfwxB
3gR+SEp+fJbQ1lRJTW84pBRrNgpgzQXiUkAkeLT0MGT9rS2L1PN9uY/fsB4qkiI3
u57pxJGmIlnLYlaqcHn9PIyI3PoG0fo4V0mDCWPEFpT2w9L5es4czqrr5Rn908pu
17sImClNtK2nYxJxuj8ZoRtZDjHauYQWXCkpwcKBeWpA57Y/hXFVdES7+TBHp+JK
jby4odzlggf7PuPnK7au1wcmSsyJTNE5lwFtnzGHDUIEJUnoTUxSGGj6OHuw9qU9
DTLMCDkBGvcSHoLdGVdvYNCxecew8qw6ee555WExABB5YzED14DCnTKyW1o/Gthp
dnFfno0RoXNZxcaSzmisAlosx0GrpQj8ReSttDKJWMHPgL3tPhUsuHUp39A4kNUc
dlQo6aEYKSlZ7cgKqeokqE9kie+KtEsVRqGZm7ys7GQv1DMpVYrswQb2hoyTw2J1
RwdMZG3Tuwh+hZjE526xW5VK7hwagCOpm5R4Xd3VN6qqsiUiusMvjU2rn8UDW2rv
t29yiUGgUt3ksrB3wK+Mofc+5Os1MGW1GXaKSTOq/p0PGbcl2djIb1+zoiEKf3mY
JJfmoNxZp0eZAPHJLvNagSG1jzGgpFYagHU2lUs5mnXBMX7PSDpc/HNm/EImUL9A
Ghb/hyaiWzSAJrsBGLseUBEkvbsJDoXHsGLI0QrjXSu1z+EatdxPrVw6mtIKHvtb
KziNY+952+hwcivyo6nZluN+OgssSU2D1lih/slBxAbICzBBVzWJMgXoI67798D4
h48bYf+mAv0Rx6ikfLnsw7dt48joqtXFAhgcMxJQ5JZeTL2g8esCh+vRINtf4cYE
MhSf0H2Ys82hmUELUq5USMojgZyWwd/5AgFC31Epq5NkvfYVWZWb4CHIODl9zfcC
hIBGWlBtXB+FdlHY1lQkBtG9+VXZPMe9HBpg1WmrNzHxlBWYPc9PncO6M7k3+2E3
V7Z3Fct67r74PJV7L7oH2EIYot+p7cyeMS9hhvrhDXneWJP7cZTN/SUTSSLe4b2u
PZYXOu6eUGwL2+00CTHjuhJL3ylPdjksfutodu+hXU1HN48oFGiS+OI+JkgR8/n4
skNc+l54TPzS3hLyDsZReUgMX3ByJmhKm/9sEywvMGkAPX/QsdMAVHBpYfb6uAwY
5WugPlYlrPTHp+Ym6nDlnsHjXhp+xusvVlLt6AFbX8ohJ8ZfjHkBT9Pufy/+uw68
PPDhMse1Zpo9gTBo/SNB71Ywl1Zv4pqOmS8B91oFzbGi0qhxeLBfjFjOLemjLD3y
8klVaai1RIQmK+ZBIZ2t9yds05ITGVza1AAu9zCBXHaGTM8KMqp3zCqCn0ddSvmw
L8H96E5Onb3fyEQ3t6PteVdIUL+1cvkn1ZJqXmNG9ZvX06HmjIo3BBKOBE3fBJkg
zXQiSAH9xvYMSKbgAo36ENwOZJ0E9DM9SQK4rdFbRt2MIx0NCtbw+Ezt92fKKhMp
PsOnx+Yinucx1qHBS5LpHQhLzd1aq7yFWt6KB2tHALsk4LEweeSxuUhMwf+BprIY
wa5cms5IZH29cEJfrizlo3EVpX4DBBaUdR5J4PINfbszcZj6dHKePITwh/Pejg7y
RUX8kv7CeifjJ59+gLMS8OjAq0EeIFmc2AHwh8CYUqxQtxe1dnA2BNNeePaLYMDn
LavOnon0ZhmXd7vjQNWWDfHwZ7ORE4JMQoLm5cSqFGjEZBre1+8xDpup/mo8k/Rw
jMgYjgAw7q51hGd5vHZSU9RF0vCdyanUyqMtRKWOeLzVWdy7++J6m/th9NsS5HaD
nDn4Bm65OssnSse3x4eiuxTOTP8S9cO52XkmphyDC4aerFeaKvMjqsNN9vBSXnHU
IYL2wA+gMpjIld7xXwegmaQPwcFL8HGBCI2kbRWSh54mKS3P2mRXOR9mc9btfTlX
H+50byHtGfbB3CpxpNEUBbvxpHoWw4P2v5idSpMnlaNlGtAeAjxwFF+RHhGzGgf0
2Q6kUhdd8bVphI542jlb1rmiyrF1LVuMUmV6SffXJVnPIA+Cz2Wyo2Y0twSl03vw
X+oxLXGIpPMsfAM6fyyiPWlN3yo6roY8fODAj2NFh9oeScUNCGnrvv3HTyz2TS7A
YTd4tK7jFwrZKvaBzy/eHbGxXeX6XRAX/noT/QD8Lm9PZQV51qlGy0fBs+oK7Lkz
l+65tL9zFO5gHtU1Xi92xoyjA5YzfMSq8OGJgv7vbzr11R4cjgCRXk+gxKN72Sho
WFrlrGoLNaVx9e/KkxNKpT2Y1VXSMgxNocAjUEGblC1mMkokbunE4tKROXFTk9Ge
G3tcmx2WPxYE3iY8BmUme8OVRI3NQ7M68I2zngyjUXjjAqtAYjD/kSDDsA9+isvv
lgmcJmbQUW9Lm9H56cicrQ==
`protect end_protected