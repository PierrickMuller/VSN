--------------------------------------------------------------------------------
-- HEIG-VD
-- Haute Ecole d'Ingenerie et de Gestion du Canton de Vaud
-- School of Business and Engineering in Canton de Vaud
--------------------------------------------------------------------------------
-- REDS Institute
-- Reconfigurable Embedded Digital Systems
--------------------------------------------------------------------------------
--
-- File     : transactions_pkg.vhd
-- Author   : Yann Thoma
-- Date     : 31.03.2021
--
-- Context  :
--
--------------------------------------------------------------------------------
-- Description : This package offers the transaction types for the Morse
--               burst emitter.
--
--------------------------------------------------------------------------------
-- Dependencies : -
--
--------------------------------------------------------------------------------
-- Modifications :
-- Ver   Date        Person     Comments
-- 0.1   31.03.2021  YTA        Initial version
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package transactions_pkg is

    -- The commands the sequencer can sends to the driver
    type command_t is (
        -- Starts a burst transmission
        send,
        -- Adds a character in the internal FIFO
        add_char,
        -- Does nothing
        nop
    );

    -- The transaction sent by the sequencer to the driver
    type input_transaction_t is record
        -- The command to be played by the driver
        command : command_t;
        -- The ASCII character to send
        char : std_logic_vector(7 downto 0);
        -- A waiting time... Maybe useful
        waiting_time : integer;
        -- A validity... Maybe useful
        valid : boolean;
        -- A dot period, used when we start a burst transmission
        dot_period : std_logic_vector(27 downto 0);
    end record;

    -- The transaction generated by the output monitor
    type output_transaction_t is record
        -- The ASCII character decoded
        char : std_logic_vector(7 downto 0);
        -- Is this character valid or not?
        valid : std_logic;
    end record;

end package;
