// Size of data, to be used everywhere
`define DATASIZE 16
